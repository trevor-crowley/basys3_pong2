`timescale 1 ns / 1 ps

module AESL_deadlock_kernel_monitor_top ( 
    input wire kernel_monitor_clock,
    input wire kernel_monitor_reset
);
wire [4:0] axis_block_sigs;
wire [13:0] inst_idle_sigs;
wire [4:0] inst_block_sigs;
wire kernel_block;

assign axis_block_sigs[0] = ~AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.grp_AXIVideo2BayerMat_0_4320_3848_2_3_Pipeline_loop_start_hunt_fu_179.in_ptr_TDATA_blk_n;
assign axis_block_sigs[1] = ~AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.grp_AXIVideo2BayerMat_0_4320_3848_2_3_Pipeline_loop_col_zxi2mat_fu_199.in_ptr_TDATA_blk_n;
assign axis_block_sigs[2] = ~AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.grp_AXIVideo2BayerMat_0_4320_3848_2_3_Pipeline_loop_last_hunt_fu_226.in_ptr_TDATA_blk_n;
assign axis_block_sigs[3] = ~AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_U0.grp_GRAYMat2AXIvideo_0_2160_3840_2_3_Pipeline_loop_col_mat2axi_fu_100.lef_ptr_TDATA_blk_n;
assign axis_block_sigs[4] = ~AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_1_U0.grp_GRAYMat2AXIvideo_0_2160_3840_2_3_1_Pipeline_loop_col_mat2axi_fu_88.sef_ptr_TDATA_blk_n;

assign inst_idle_sigs[0] = AESL_inst_extractEFrames_accel.Block_entry5_proc_U0.ap_idle;
assign inst_block_sigs[0] = (AESL_inst_extractEFrames_accel.Block_entry5_proc_U0.ap_done & ~AESL_inst_extractEFrames_accel.Block_entry5_proc_U0.ap_continue);
assign inst_idle_sigs[1] = AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.ap_idle;
assign inst_block_sigs[1] = (AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.ap_done & ~AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.ap_continue) | ~AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.grp_AXIVideo2BayerMat_0_4320_3848_2_3_Pipeline_loop_col_zxi2mat_fu_199.InImg_data156_blk_n | ~AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.InImg_cols_c_blk_n;
assign inst_idle_sigs[2] = AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.ap_idle;
assign inst_block_sigs[2] = (AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.ap_done & ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.ap_continue) | ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.p_hdrSrc_cols_blk_n | ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.grp_extract_fu_102.grp_extract_Pipeline_LAST_LINES_VITIS_LOOP_177_4_fu_190.InImg_data156_blk_n | ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.grp_extract_fu_102.grp_extract_Pipeline_VITIS_LOOP_145_3_fu_162.InImg_data156_blk_n | ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.grp_extract_fu_102.grp_extract_Pipeline_VITIS_LOOP_133_2_fu_138.InImg_data156_blk_n | ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.grp_extract_fu_102.grp_extract_Pipeline_VITIS_LOOP_113_1_fu_116.InImg_data156_blk_n | ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.grp_extract_fu_102.grp_extract_Pipeline_LAST_LINES_VITIS_LOOP_177_4_fu_190.LEF_Img_data157_blk_n | ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.grp_extract_fu_102.grp_extract_Pipeline_VITIS_LOOP_145_3_fu_162.LEF_Img_data157_blk_n | ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.grp_extract_fu_102.grp_extract_Pipeline_LAST_LINES_VITIS_LOOP_177_4_fu_190.SEF_Img_data158_blk_n | ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.grp_extract_fu_102.grp_extract_Pipeline_VITIS_LOOP_145_3_fu_162.SEF_Img_data158_blk_n | ~AESL_inst_extractEFrames_accel.extractExposureFrames_0_8_8_2160_3840_2_3_3_3_0_U0.LEF_Img_rows_c_blk_n;
assign inst_idle_sigs[3] = AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_U0.ap_idle;
assign inst_block_sigs[3] = (AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_U0.ap_done & ~AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_U0.ap_continue) | ~AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_U0.gray_mat_rows_blk_n | ~AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_U0.grp_GRAYMat2AXIvideo_0_2160_3840_2_3_Pipeline_loop_col_mat2axi_fu_100.LEF_Img_data157_blk_n;
assign inst_idle_sigs[4] = AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_1_U0.ap_idle;
assign inst_block_sigs[4] = (AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_1_U0.ap_done & ~AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_1_U0.ap_continue) | ~AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_1_U0.grp_GRAYMat2AXIvideo_0_2160_3840_2_3_1_Pipeline_loop_col_mat2axi_fu_88.SEF_Img_data158_blk_n;

assign inst_idle_sigs[5] = 1'b0;
assign inst_idle_sigs[6] = AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.ap_idle;
assign inst_idle_sigs[7] = AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.grp_AXIVideo2BayerMat_0_4320_3848_2_3_Pipeline_loop_start_hunt_fu_179.ap_idle;
assign inst_idle_sigs[8] = AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.grp_AXIVideo2BayerMat_0_4320_3848_2_3_Pipeline_loop_col_zxi2mat_fu_199.ap_idle;
assign inst_idle_sigs[9] = AESL_inst_extractEFrames_accel.AXIVideo2BayerMat_0_4320_3848_2_3_U0.grp_AXIVideo2BayerMat_0_4320_3848_2_3_Pipeline_loop_last_hunt_fu_226.ap_idle;
assign inst_idle_sigs[10] = AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_U0.ap_idle;
assign inst_idle_sigs[11] = AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_U0.grp_GRAYMat2AXIvideo_0_2160_3840_2_3_Pipeline_loop_col_mat2axi_fu_100.ap_idle;
assign inst_idle_sigs[12] = AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_1_U0.ap_idle;
assign inst_idle_sigs[13] = AESL_inst_extractEFrames_accel.GRAYMat2AXIvideo_0_2160_3840_2_3_1_U0.grp_GRAYMat2AXIvideo_0_2160_3840_2_3_1_Pipeline_loop_col_mat2axi_fu_88.ap_idle;

AESL_deadlock_idx0_monitor AESL_deadlock_idx0_monitor_U (
    .clock(kernel_monitor_clock),
    .reset(kernel_monitor_reset),
    .axis_block_sigs(axis_block_sigs),
    .inst_idle_sigs(inst_idle_sigs),
    .inst_block_sigs(inst_block_sigs),
    .block(kernel_block)
);

initial begin
reg block_delay = 0;
    while(1) begin
        @(posedge kernel_monitor_clock);
    if (kernel_block == 1'b1 && block_delay == 1'b0)
    $display("find kernel block.");
    block_delay = kernel_block;
    end
end

endmodule
